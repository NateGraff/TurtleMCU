
module rom(
	input wire [9:0] addr,
	output wire [15:0] dout);

	assign dout = 16'h0000;

endmodule